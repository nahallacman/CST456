`timescale 1 ns / 1 ns // timescale for following modules

// Change MAX_INDEX to 256 for your program.
`define MAX_INDEX 256

// The RAM block that stores the program to be run by the 68HC11.
module int_ram
(
	E,
	rw,
	address,
	data_in,
	data_out
);

	input E;
	input rw;
	input [15:0] address;
	input [7:0] data_in;
	output [7:0] data_out;

	reg [7:0] ram[65535:0];
	
	// Put program here. This is the output of your conversion script.
	initial
	begin
ram[8192] = 8'h86;
ram[8193] = 8'h00;
ram[8194] = 8'h43;
ram[8195] = 8'hB7;
ram[8196] = 8'h40;
ram[8197] = 8'h00;
ram[8198] = 8'h86;
ram[8199] = 8'h01;
ram[8200] = 8'h43;
ram[8201] = 8'hB7;
ram[8202] = 8'h40;
ram[8203] = 8'h01;
ram[8204] = 8'h86;
ram[8205] = 8'h02;
ram[8206] = 8'h43;
ram[8207] = 8'hB7;
ram[8208] = 8'h40;
ram[8209] = 8'h02;
ram[8210] = 8'h86;
ram[8211] = 8'h03;
ram[8212] = 8'h43;
ram[8213] = 8'hB7;
ram[8214] = 8'h40;
ram[8215] = 8'h03;
ram[8216] = 8'h86;
ram[8217] = 8'h04;
ram[8218] = 8'h43;
ram[8219] = 8'hB7;
ram[8220] = 8'h40;
ram[8221] = 8'h04;
ram[8222] = 8'h86;
ram[8223] = 8'h05;
ram[8224] = 8'h43;
ram[8225] = 8'hB7;
ram[8226] = 8'h40;
ram[8227] = 8'h05;
ram[8228] = 8'h86;
ram[8229] = 8'h06;
ram[8230] = 8'h43;
ram[8231] = 8'hB7;
ram[8232] = 8'h40;
ram[8233] = 8'h06;
ram[8234] = 8'h86;
ram[8235] = 8'h07;
ram[8236] = 8'h43;
ram[8237] = 8'hB7;
ram[8238] = 8'h40;
ram[8239] = 8'h07;
ram[8240] = 8'h86;
ram[8241] = 8'h08;
ram[8242] = 8'h43;
ram[8243] = 8'hB7;
ram[8244] = 8'h40;
ram[8245] = 8'h08;
ram[8246] = 8'h86;
ram[8247] = 8'h09;
ram[8248] = 8'h43;
ram[8249] = 8'hB7;
ram[8250] = 8'h40;
ram[8251] = 8'h09;
ram[8252] = 8'h86;
ram[8253] = 8'h0A;
ram[8254] = 8'h43;
ram[8255] = 8'hB7;
ram[8256] = 8'h40;
ram[8257] = 8'h0A;
ram[8258] = 8'h86;
ram[8259] = 8'h0B;
ram[8260] = 8'h43;
ram[8261] = 8'hB7;
ram[8262] = 8'h40;
ram[8263] = 8'h0B;
ram[8264] = 8'h86;
ram[8265] = 8'h0C;
ram[8266] = 8'h43;
ram[8267] = 8'hB7;
ram[8268] = 8'h40;
ram[8269] = 8'h0C;
ram[8270] = 8'h86;
ram[8271] = 8'h0D;
ram[8272] = 8'h43;
ram[8273] = 8'hB7;
ram[8274] = 8'h40;
ram[8275] = 8'h0D;
ram[8276] = 8'h86;
ram[8277] = 8'h0E;
ram[8278] = 8'h43;
ram[8279] = 8'hB7;
ram[8280] = 8'h40;
ram[8281] = 8'h0E;
ram[8282] = 8'h86;
ram[8283] = 8'h0F;
ram[8284] = 8'h43;
ram[8285] = 8'hB7;
ram[8286] = 8'h40;
ram[8287] = 8'h0F;
ram[8288] = 8'h86;
ram[8289] = 8'h10;
ram[8290] = 8'h43;
ram[8291] = 8'hB7;
ram[8292] = 8'h40;
ram[8293] = 8'h10;
ram[8294] = 8'h86;
ram[8295] = 8'h11;
ram[8296] = 8'h43;
ram[8297] = 8'hB7;
ram[8298] = 8'h40;
ram[8299] = 8'h11;
ram[8300] = 8'h86;
ram[8301] = 8'h12;
ram[8302] = 8'h43;
ram[8303] = 8'hB7;
ram[8304] = 8'h40;
ram[8305] = 8'h12;
ram[8306] = 8'h86;
ram[8307] = 8'h13;
ram[8308] = 8'h43;
ram[8309] = 8'hB7;
ram[8310] = 8'h40;
ram[8311] = 8'h13;
ram[8312] = 8'h86;
ram[8313] = 8'h14;
ram[8314] = 8'h43;
ram[8315] = 8'hB7;
ram[8316] = 8'h40;
ram[8317] = 8'h14;
ram[8318] = 8'h86;
ram[8319] = 8'h15;
ram[8320] = 8'h43;
ram[8321] = 8'hB7;
ram[8322] = 8'h40;
ram[8323] = 8'h15;
ram[8324] = 8'h86;
ram[8325] = 8'h16;
ram[8326] = 8'h43;
ram[8327] = 8'hB7;
ram[8328] = 8'h40;
ram[8329] = 8'h16;
ram[8330] = 8'h86;
ram[8331] = 8'h17;
ram[8332] = 8'h43;
ram[8333] = 8'hB7;
ram[8334] = 8'h40;
ram[8335] = 8'h17;
ram[8336] = 8'h86;
ram[8337] = 8'h18;
ram[8338] = 8'h43;
ram[8339] = 8'hB7;
ram[8340] = 8'h40;
ram[8341] = 8'h18;
ram[8342] = 8'h86;
ram[8343] = 8'h19;
ram[8344] = 8'h43;
ram[8345] = 8'hB7;
ram[8346] = 8'h40;
ram[8347] = 8'h19;
ram[8348] = 8'h86;
ram[8349] = 8'h1A;
ram[8350] = 8'h43;
ram[8351] = 8'hB7;
ram[8352] = 8'h40;
ram[8353] = 8'h1A;
ram[8354] = 8'h86;
ram[8355] = 8'h1B;
ram[8356] = 8'h43;
ram[8357] = 8'hB7;
ram[8358] = 8'h40;
ram[8359] = 8'h1B;
ram[8360] = 8'h86;
ram[8361] = 8'h1C;
ram[8362] = 8'h43;
ram[8363] = 8'hB7;
ram[8364] = 8'h40;
ram[8365] = 8'h1C;
ram[8366] = 8'h86;
ram[8367] = 8'h1D;
ram[8368] = 8'h43;
ram[8369] = 8'hB7;
ram[8370] = 8'h40;
ram[8371] = 8'h1D;
ram[8372] = 8'h86;
ram[8373] = 8'h1E;
ram[8374] = 8'h43;
ram[8375] = 8'hB7;
ram[8376] = 8'h40;
ram[8377] = 8'h1E;
ram[8378] = 8'h86;
ram[8379] = 8'h1F;
ram[8380] = 8'h43;
ram[8381] = 8'hB7;
ram[8382] = 8'h40;
ram[8383] = 8'h1F;
ram[8384] = 8'h86;
ram[8385] = 8'h20;
ram[8386] = 8'h43;
ram[8387] = 8'hB7;
ram[8388] = 8'h40;
ram[8389] = 8'h20;
ram[8390] = 8'h86;
ram[8391] = 8'h21;
ram[8392] = 8'h43;
ram[8393] = 8'hB7;
ram[8394] = 8'h40;
ram[8395] = 8'h21;
ram[8396] = 8'h86;
ram[8397] = 8'h22;
ram[8398] = 8'h43;
ram[8399] = 8'hB7;
ram[8400] = 8'h40;
ram[8401] = 8'h22;
ram[8402] = 8'h86;
ram[8403] = 8'h23;
ram[8404] = 8'h43;
ram[8405] = 8'hB7;
ram[8406] = 8'h40;
ram[8407] = 8'h23;
ram[8408] = 8'h86;
ram[8409] = 8'h24;
ram[8410] = 8'h43;
ram[8411] = 8'hB7;
ram[8412] = 8'h40;
ram[8413] = 8'h24;
ram[8414] = 8'h86;
ram[8415] = 8'h25;
ram[8416] = 8'h43;
ram[8417] = 8'hB7;
ram[8418] = 8'h40;
ram[8419] = 8'h25;
ram[8420] = 8'h86;
ram[8421] = 8'h26;
ram[8422] = 8'h43;
ram[8423] = 8'hB7;
ram[8424] = 8'h40;
ram[8425] = 8'h26;
ram[8426] = 8'h86;
ram[8427] = 8'h27;
ram[8428] = 8'h43;
ram[8429] = 8'hB7;
ram[8430] = 8'h40;
ram[8431] = 8'h27;
ram[8432] = 8'h86;
ram[8433] = 8'h28;
ram[8434] = 8'h43;
ram[8435] = 8'hB7;
ram[8436] = 8'h40;
ram[8437] = 8'h28;
ram[8438] = 8'h86;
ram[8439] = 8'h29;
ram[8440] = 8'h43;
ram[8441] = 8'hB7;
ram[8442] = 8'h40;
ram[8443] = 8'h29;
ram[8444] = 8'h86;
ram[8445] = 8'h2A;
ram[8446] = 8'h43;
ram[8447] = 8'hB7;
ram[8448] = 8'h40;
ram[8449] = 8'h2A;
ram[8450] = 8'h86;
ram[8451] = 8'h2B;
ram[8452] = 8'h43;
ram[8453] = 8'hB7;
ram[8454] = 8'h40;
ram[8455] = 8'h2B;
ram[8456] = 8'h86;
ram[8457] = 8'h2C;
ram[8458] = 8'h43;
ram[8459] = 8'hB7;
ram[8460] = 8'h40;
ram[8461] = 8'h2C;
ram[8462] = 8'h86;
ram[8463] = 8'h2D;
ram[8464] = 8'h43;
ram[8465] = 8'hB7;
ram[8466] = 8'h40;
ram[8467] = 8'h2D;
ram[8468] = 8'h86;
ram[8469] = 8'h2E;
ram[8470] = 8'h43;
ram[8471] = 8'hB7;
ram[8472] = 8'h40;
ram[8473] = 8'h2E;
ram[8474] = 8'h86;
ram[8475] = 8'h2F;
ram[8476] = 8'h43;
ram[8477] = 8'hB7;
ram[8478] = 8'h40;
ram[8479] = 8'h2F;
ram[8480] = 8'h86;
ram[8481] = 8'h30;
ram[8482] = 8'h43;
ram[8483] = 8'hB7;
ram[8484] = 8'h40;
ram[8485] = 8'h30;
ram[8486] = 8'h86;
ram[8487] = 8'h31;
ram[8488] = 8'h43;
ram[8489] = 8'hB7;
ram[8490] = 8'h40;
ram[8491] = 8'h31;
ram[8492] = 8'h86;
ram[8493] = 8'h32;
ram[8494] = 8'h43;
ram[8495] = 8'hB7;
ram[8496] = 8'h40;
ram[8497] = 8'h32;
ram[8498] = 8'h86;
ram[8499] = 8'h33;
ram[8500] = 8'h43;
ram[8501] = 8'hB7;
ram[8502] = 8'h40;
ram[8503] = 8'h33;
ram[8504] = 8'h86;
ram[8505] = 8'h34;
ram[8506] = 8'h43;
ram[8507] = 8'hB7;
ram[8508] = 8'h40;
ram[8509] = 8'h34;
ram[8510] = 8'h86;
ram[8511] = 8'h35;
ram[8512] = 8'h43;
ram[8513] = 8'hB7;
ram[8514] = 8'h40;
ram[8515] = 8'h35;
ram[8516] = 8'h86;
ram[8517] = 8'h36;
ram[8518] = 8'h43;
ram[8519] = 8'hB7;
ram[8520] = 8'h40;
ram[8521] = 8'h36;
ram[8522] = 8'h86;
ram[8523] = 8'h37;
ram[8524] = 8'h43;
ram[8525] = 8'hB7;
ram[8526] = 8'h40;
ram[8527] = 8'h37;
ram[8528] = 8'h86;
ram[8529] = 8'h38;
ram[8530] = 8'h43;
ram[8531] = 8'hB7;
ram[8532] = 8'h40;
ram[8533] = 8'h38;
ram[8534] = 8'h86;
ram[8535] = 8'h39;
ram[8536] = 8'h43;
ram[8537] = 8'hB7;
ram[8538] = 8'h40;
ram[8539] = 8'h39;
ram[8540] = 8'h86;
ram[8541] = 8'h3A;
ram[8542] = 8'h43;
ram[8543] = 8'hB7;
ram[8544] = 8'h40;
ram[8545] = 8'h3A;
ram[8546] = 8'h86;
ram[8547] = 8'h3B;
ram[8548] = 8'h43;
ram[8549] = 8'hB7;
ram[8550] = 8'h40;
ram[8551] = 8'h3B;
ram[8552] = 8'h86;
ram[8553] = 8'h3C;
ram[8554] = 8'h43;
ram[8555] = 8'hB7;
ram[8556] = 8'h40;
ram[8557] = 8'h3C;
ram[8558] = 8'h86;
ram[8559] = 8'h3D;
ram[8560] = 8'h43;
ram[8561] = 8'hB7;
ram[8562] = 8'h40;
ram[8563] = 8'h3D;
ram[8564] = 8'h86;
ram[8565] = 8'h3E;
ram[8566] = 8'h43;
ram[8567] = 8'hB7;
ram[8568] = 8'h40;
ram[8569] = 8'h3E;
ram[8570] = 8'h86;
ram[8571] = 8'h3F;
ram[8572] = 8'h43;
ram[8573] = 8'hB7;
ram[8574] = 8'h40;
ram[8575] = 8'h3F;
ram[8576] = 8'h86;
ram[8577] = 8'h40;
ram[8578] = 8'h43;
ram[8579] = 8'hB7;
ram[8580] = 8'h40;
ram[8581] = 8'h40;
ram[8582] = 8'h86;
ram[8583] = 8'h41;
ram[8584] = 8'h43;
ram[8585] = 8'hB7;
ram[8586] = 8'h40;
ram[8587] = 8'h41;
ram[8588] = 8'h86;
ram[8589] = 8'h42;
ram[8590] = 8'h43;
ram[8591] = 8'hB7;
ram[8592] = 8'h40;
ram[8593] = 8'h42;
ram[8594] = 8'h86;
ram[8595] = 8'h43;
ram[8596] = 8'h43;
ram[8597] = 8'hB7;
ram[8598] = 8'h40;
ram[8599] = 8'h43;
ram[8600] = 8'h86;
ram[8601] = 8'h44;
ram[8602] = 8'h43;
ram[8603] = 8'hB7;
ram[8604] = 8'h40;
ram[8605] = 8'h44;
ram[8606] = 8'h86;
ram[8607] = 8'h45;
ram[8608] = 8'h43;
ram[8609] = 8'hB7;
ram[8610] = 8'h40;
ram[8611] = 8'h45;
ram[8612] = 8'h86;
ram[8613] = 8'h46;
ram[8614] = 8'h43;
ram[8615] = 8'hB7;
ram[8616] = 8'h40;
ram[8617] = 8'h46;
ram[8618] = 8'h86;
ram[8619] = 8'h47;
ram[8620] = 8'h43;
ram[8621] = 8'hB7;
ram[8622] = 8'h40;
ram[8623] = 8'h47;
ram[8624] = 8'h86;
ram[8625] = 8'h48;
ram[8626] = 8'h43;
ram[8627] = 8'hB7;
ram[8628] = 8'h40;
ram[8629] = 8'h48;
ram[8630] = 8'h86;
ram[8631] = 8'h49;
ram[8632] = 8'h43;
ram[8633] = 8'hB7;
ram[8634] = 8'h40;
ram[8635] = 8'h49;
ram[8636] = 8'h86;
ram[8637] = 8'h4A;
ram[8638] = 8'h43;
ram[8639] = 8'hB7;
ram[8640] = 8'h40;
ram[8641] = 8'h4A;
ram[8642] = 8'h86;
ram[8643] = 8'h4B;
ram[8644] = 8'h43;
ram[8645] = 8'hB7;
ram[8646] = 8'h40;
ram[8647] = 8'h4B;
ram[8648] = 8'h86;
ram[8649] = 8'h4C;
ram[8650] = 8'h43;
ram[8651] = 8'hB7;
ram[8652] = 8'h40;
ram[8653] = 8'h4C;
ram[8654] = 8'h86;
ram[8655] = 8'h4D;
ram[8656] = 8'h43;
ram[8657] = 8'hB7;
ram[8658] = 8'h40;
ram[8659] = 8'h4D;
ram[8660] = 8'h86;
ram[8661] = 8'h4E;
ram[8662] = 8'h43;
ram[8663] = 8'hB7;
ram[8664] = 8'h40;
ram[8665] = 8'h4E;
ram[8666] = 8'h86;
ram[8667] = 8'h4F;
ram[8668] = 8'h43;
ram[8669] = 8'hB7;
ram[8670] = 8'h40;
ram[8671] = 8'h4F;
ram[8672] = 8'h86;
ram[8673] = 8'h50;
ram[8674] = 8'h43;
ram[8675] = 8'hB7;
ram[8676] = 8'h40;
ram[8677] = 8'h50;
ram[8678] = 8'h86;
ram[8679] = 8'h51;
ram[8680] = 8'h43;
ram[8681] = 8'hB7;
ram[8682] = 8'h40;
ram[8683] = 8'h51;
ram[8684] = 8'h86;
ram[8685] = 8'h52;
ram[8686] = 8'h43;
ram[8687] = 8'hB7;
ram[8688] = 8'h40;
ram[8689] = 8'h52;
ram[8690] = 8'h86;
ram[8691] = 8'h53;
ram[8692] = 8'h43;
ram[8693] = 8'hB7;
ram[8694] = 8'h40;
ram[8695] = 8'h53;
ram[8696] = 8'h86;
ram[8697] = 8'h54;
ram[8698] = 8'h43;
ram[8699] = 8'hB7;
ram[8700] = 8'h40;
ram[8701] = 8'h54;
ram[8702] = 8'h86;
ram[8703] = 8'h55;
ram[8704] = 8'h43;
ram[8705] = 8'hB7;
ram[8706] = 8'h40;
ram[8707] = 8'h55;
ram[8708] = 8'h86;
ram[8709] = 8'h56;
ram[8710] = 8'h43;
ram[8711] = 8'hB7;
ram[8712] = 8'h40;
ram[8713] = 8'h56;
ram[8714] = 8'h86;
ram[8715] = 8'h57;
ram[8716] = 8'h43;
ram[8717] = 8'hB7;
ram[8718] = 8'h40;
ram[8719] = 8'h57;
ram[8720] = 8'h86;
ram[8721] = 8'h58;
ram[8722] = 8'h43;
ram[8723] = 8'hB7;
ram[8724] = 8'h40;
ram[8725] = 8'h58;
ram[8726] = 8'h86;
ram[8727] = 8'h59;
ram[8728] = 8'h43;
ram[8729] = 8'hB7;
ram[8730] = 8'h40;
ram[8731] = 8'h59;
ram[8732] = 8'h86;
ram[8733] = 8'h5A;
ram[8734] = 8'h43;
ram[8735] = 8'hB7;
ram[8736] = 8'h40;
ram[8737] = 8'h5A;
ram[8738] = 8'h86;
ram[8739] = 8'h5B;
ram[8740] = 8'h43;
ram[8741] = 8'hB7;
ram[8742] = 8'h40;
ram[8743] = 8'h5B;
ram[8744] = 8'h86;
ram[8745] = 8'h5C;
ram[8746] = 8'h43;
ram[8747] = 8'hB7;
ram[8748] = 8'h40;
ram[8749] = 8'h5C;
ram[8750] = 8'h86;
ram[8751] = 8'h5D;
ram[8752] = 8'h43;
ram[8753] = 8'hB7;
ram[8754] = 8'h40;
ram[8755] = 8'h5D;
ram[8756] = 8'h86;
ram[8757] = 8'h5E;
ram[8758] = 8'h43;
ram[8759] = 8'hB7;
ram[8760] = 8'h40;
ram[8761] = 8'h5E;
ram[8762] = 8'h86;
ram[8763] = 8'h5F;
ram[8764] = 8'h43;
ram[8765] = 8'hB7;
ram[8766] = 8'h40;
ram[8767] = 8'h5F;
ram[8768] = 8'h86;
ram[8769] = 8'h60;
ram[8770] = 8'h43;
ram[8771] = 8'hB7;
ram[8772] = 8'h40;
ram[8773] = 8'h60;
ram[8774] = 8'h86;
ram[8775] = 8'h61;
ram[8776] = 8'h43;
ram[8777] = 8'hB7;
ram[8778] = 8'h40;
ram[8779] = 8'h61;
ram[8780] = 8'h86;
ram[8781] = 8'h62;
ram[8782] = 8'h43;
ram[8783] = 8'hB7;
ram[8784] = 8'h40;
ram[8785] = 8'h62;
ram[8786] = 8'h86;
ram[8787] = 8'h63;
ram[8788] = 8'h43;
ram[8789] = 8'hB7;
ram[8790] = 8'h40;
ram[8791] = 8'h63;
ram[8792] = 8'h86;
ram[8793] = 8'h64;
ram[8794] = 8'h43;
ram[8795] = 8'hB7;
ram[8796] = 8'h40;
ram[8797] = 8'h64;
ram[8798] = 8'h86;
ram[8799] = 8'h65;
ram[8800] = 8'h43;
ram[8801] = 8'hB7;
ram[8802] = 8'h40;
ram[8803] = 8'h65;
ram[8804] = 8'h86;
ram[8805] = 8'h66;
ram[8806] = 8'h43;
ram[8807] = 8'hB7;
ram[8808] = 8'h40;
ram[8809] = 8'h66;
ram[8810] = 8'h86;
ram[8811] = 8'h67;
ram[8812] = 8'h43;
ram[8813] = 8'hB7;
ram[8814] = 8'h40;
ram[8815] = 8'h67;
ram[8816] = 8'h86;
ram[8817] = 8'h68;
ram[8818] = 8'h43;
ram[8819] = 8'hB7;
ram[8820] = 8'h40;
ram[8821] = 8'h68;
ram[8822] = 8'h86;
ram[8823] = 8'h69;
ram[8824] = 8'h43;
ram[8825] = 8'hB7;
ram[8826] = 8'h40;
ram[8827] = 8'h69;
ram[8828] = 8'h86;
ram[8829] = 8'h6A;
ram[8830] = 8'h43;
ram[8831] = 8'hB7;
ram[8832] = 8'h40;
ram[8833] = 8'h6A;
ram[8834] = 8'h86;
ram[8835] = 8'h6B;
ram[8836] = 8'h43;
ram[8837] = 8'hB7;
ram[8838] = 8'h40;
ram[8839] = 8'h6B;
ram[8840] = 8'h86;
ram[8841] = 8'h6C;
ram[8842] = 8'h43;
ram[8843] = 8'hB7;
ram[8844] = 8'h40;
ram[8845] = 8'h6C;
ram[8846] = 8'h86;
ram[8847] = 8'h6D;
ram[8848] = 8'h43;
ram[8849] = 8'hB7;
ram[8850] = 8'h40;
ram[8851] = 8'h6D;
ram[8852] = 8'h86;
ram[8853] = 8'h6E;
ram[8854] = 8'h43;
ram[8855] = 8'hB7;
ram[8856] = 8'h40;
ram[8857] = 8'h6E;
ram[8858] = 8'h86;
ram[8859] = 8'h6F;
ram[8860] = 8'h43;
ram[8861] = 8'hB7;
ram[8862] = 8'h40;
ram[8863] = 8'h6F;
ram[8864] = 8'h86;
ram[8865] = 8'h70;
ram[8866] = 8'h43;
ram[8867] = 8'hB7;
ram[8868] = 8'h40;
ram[8869] = 8'h70;
ram[8870] = 8'h86;
ram[8871] = 8'h71;
ram[8872] = 8'h43;
ram[8873] = 8'hB7;
ram[8874] = 8'h40;
ram[8875] = 8'h71;
ram[8876] = 8'h86;
ram[8877] = 8'h72;
ram[8878] = 8'h43;
ram[8879] = 8'hB7;
ram[8880] = 8'h40;
ram[8881] = 8'h72;
ram[8882] = 8'h86;
ram[8883] = 8'h73;
ram[8884] = 8'h43;
ram[8885] = 8'hB7;
ram[8886] = 8'h40;
ram[8887] = 8'h73;
ram[8888] = 8'h86;
ram[8889] = 8'h74;
ram[8890] = 8'h43;
ram[8891] = 8'hB7;
ram[8892] = 8'h40;
ram[8893] = 8'h74;
ram[8894] = 8'h86;
ram[8895] = 8'h75;
ram[8896] = 8'h43;
ram[8897] = 8'hB7;
ram[8898] = 8'h40;
ram[8899] = 8'h75;
ram[8900] = 8'h86;
ram[8901] = 8'h76;
ram[8902] = 8'h43;
ram[8903] = 8'hB7;
ram[8904] = 8'h40;
ram[8905] = 8'h76;
ram[8906] = 8'h86;
ram[8907] = 8'h77;
ram[8908] = 8'h43;
ram[8909] = 8'hB7;
ram[8910] = 8'h40;
ram[8911] = 8'h77;
ram[8912] = 8'h86;
ram[8913] = 8'h78;
ram[8914] = 8'h43;
ram[8915] = 8'hB7;
ram[8916] = 8'h40;
ram[8917] = 8'h78;
ram[8918] = 8'h86;
ram[8919] = 8'h79;
ram[8920] = 8'h43;
ram[8921] = 8'hB7;
ram[8922] = 8'h40;
ram[8923] = 8'h79;
ram[8924] = 8'h86;
ram[8925] = 8'h7A;
ram[8926] = 8'h43;
ram[8927] = 8'hB7;
ram[8928] = 8'h40;
ram[8929] = 8'h7A;
ram[8930] = 8'h86;
ram[8931] = 8'h7B;
ram[8932] = 8'h43;
ram[8933] = 8'hB7;
ram[8934] = 8'h40;
ram[8935] = 8'h7B;
ram[8936] = 8'h86;
ram[8937] = 8'h7C;
ram[8938] = 8'h43;
ram[8939] = 8'hB7;
ram[8940] = 8'h40;
ram[8941] = 8'h7C;
ram[8942] = 8'h86;
ram[8943] = 8'h7D;
ram[8944] = 8'h43;
ram[8945] = 8'hB7;
ram[8946] = 8'h40;
ram[8947] = 8'h7D;
ram[8948] = 8'h86;
ram[8949] = 8'h7E;
ram[8950] = 8'h43;
ram[8951] = 8'hB7;
ram[8952] = 8'h40;
ram[8953] = 8'h7E;
ram[8954] = 8'h86;
ram[8955] = 8'h7F;
ram[8956] = 8'h43;
ram[8957] = 8'hB7;
ram[8958] = 8'h40;
ram[8959] = 8'h7F;
ram[8960] = 8'h86;
ram[8961] = 8'h80;
ram[8962] = 8'h43;
ram[8963] = 8'hB7;
ram[8964] = 8'h40;
ram[8965] = 8'h80;
ram[8966] = 8'h86;
ram[8967] = 8'h81;
ram[8968] = 8'h43;
ram[8969] = 8'hB7;
ram[8970] = 8'h40;
ram[8971] = 8'h81;
ram[8972] = 8'h86;
ram[8973] = 8'h82;
ram[8974] = 8'h43;
ram[8975] = 8'hB7;
ram[8976] = 8'h40;
ram[8977] = 8'h82;
ram[8978] = 8'h86;
ram[8979] = 8'h83;
ram[8980] = 8'h43;
ram[8981] = 8'hB7;
ram[8982] = 8'h40;
ram[8983] = 8'h83;
ram[8984] = 8'h86;
ram[8985] = 8'h84;
ram[8986] = 8'h43;
ram[8987] = 8'hB7;
ram[8988] = 8'h40;
ram[8989] = 8'h84;
ram[8990] = 8'h86;
ram[8991] = 8'h85;
ram[8992] = 8'h43;
ram[8993] = 8'hB7;
ram[8994] = 8'h40;
ram[8995] = 8'h85;
ram[8996] = 8'h86;
ram[8997] = 8'h86;
ram[8998] = 8'h43;
ram[8999] = 8'hB7;
ram[9000] = 8'h40;
ram[9001] = 8'h86;
ram[9002] = 8'h86;
ram[9003] = 8'h87;
ram[9004] = 8'h43;
ram[9005] = 8'hB7;
ram[9006] = 8'h40;
ram[9007] = 8'h87;
ram[9008] = 8'h86;
ram[9009] = 8'h88;
ram[9010] = 8'h43;
ram[9011] = 8'hB7;
ram[9012] = 8'h40;
ram[9013] = 8'h88;
ram[9014] = 8'h86;
ram[9015] = 8'h89;
ram[9016] = 8'h43;
ram[9017] = 8'hB7;
ram[9018] = 8'h40;
ram[9019] = 8'h89;
ram[9020] = 8'h86;
ram[9021] = 8'h8A;
ram[9022] = 8'h43;
ram[9023] = 8'hB7;
ram[9024] = 8'h40;
ram[9025] = 8'h8A;
ram[9026] = 8'h86;
ram[9027] = 8'h8B;
ram[9028] = 8'h43;
ram[9029] = 8'hB7;
ram[9030] = 8'h40;
ram[9031] = 8'h8B;
ram[9032] = 8'h86;
ram[9033] = 8'h8C;
ram[9034] = 8'h43;
ram[9035] = 8'hB7;
ram[9036] = 8'h40;
ram[9037] = 8'h8C;
ram[9038] = 8'h86;
ram[9039] = 8'h8D;
ram[9040] = 8'h43;
ram[9041] = 8'hB7;
ram[9042] = 8'h40;
ram[9043] = 8'h8D;
ram[9044] = 8'h86;
ram[9045] = 8'h8E;
ram[9046] = 8'h43;
ram[9047] = 8'hB7;
ram[9048] = 8'h40;
ram[9049] = 8'h8E;
ram[9050] = 8'h86;
ram[9051] = 8'h8F;
ram[9052] = 8'h43;
ram[9053] = 8'hB7;
ram[9054] = 8'h40;
ram[9055] = 8'h8F;
ram[9056] = 8'h86;
ram[9057] = 8'h90;
ram[9058] = 8'h43;
ram[9059] = 8'hB7;
ram[9060] = 8'h40;
ram[9061] = 8'h90;
ram[9062] = 8'h86;
ram[9063] = 8'h91;
ram[9064] = 8'h43;
ram[9065] = 8'hB7;
ram[9066] = 8'h40;
ram[9067] = 8'h91;
ram[9068] = 8'h86;
ram[9069] = 8'h92;
ram[9070] = 8'h43;
ram[9071] = 8'hB7;
ram[9072] = 8'h40;
ram[9073] = 8'h92;
ram[9074] = 8'h86;
ram[9075] = 8'h93;
ram[9076] = 8'h43;
ram[9077] = 8'hB7;
ram[9078] = 8'h40;
ram[9079] = 8'h93;
ram[9080] = 8'h86;
ram[9081] = 8'h94;
ram[9082] = 8'h43;
ram[9083] = 8'hB7;
ram[9084] = 8'h40;
ram[9085] = 8'h94;
ram[9086] = 8'h86;
ram[9087] = 8'h95;
ram[9088] = 8'h43;
ram[9089] = 8'hB7;
ram[9090] = 8'h40;
ram[9091] = 8'h95;
ram[9092] = 8'h86;
ram[9093] = 8'h96;
ram[9094] = 8'h43;
ram[9095] = 8'hB7;
ram[9096] = 8'h40;
ram[9097] = 8'h96;
ram[9098] = 8'h86;
ram[9099] = 8'h97;
ram[9100] = 8'h43;
ram[9101] = 8'hB7;
ram[9102] = 8'h40;
ram[9103] = 8'h97;
ram[9104] = 8'h86;
ram[9105] = 8'h98;
ram[9106] = 8'h43;
ram[9107] = 8'hB7;
ram[9108] = 8'h40;
ram[9109] = 8'h98;
ram[9110] = 8'h86;
ram[9111] = 8'h99;
ram[9112] = 8'h43;
ram[9113] = 8'hB7;
ram[9114] = 8'h40;
ram[9115] = 8'h99;
ram[9116] = 8'h86;
ram[9117] = 8'h9A;
ram[9118] = 8'h43;
ram[9119] = 8'hB7;
ram[9120] = 8'h40;
ram[9121] = 8'h9A;
ram[9122] = 8'h86;
ram[9123] = 8'h9B;
ram[9124] = 8'h43;
ram[9125] = 8'hB7;
ram[9126] = 8'h40;
ram[9127] = 8'h9B;
ram[9128] = 8'h86;
ram[9129] = 8'h9C;
ram[9130] = 8'h43;
ram[9131] = 8'hB7;
ram[9132] = 8'h40;
ram[9133] = 8'h9C;
ram[9134] = 8'h86;
ram[9135] = 8'h9D;
ram[9136] = 8'h43;
ram[9137] = 8'hB7;
ram[9138] = 8'h40;
ram[9139] = 8'h9D;
ram[9140] = 8'h86;
ram[9141] = 8'h9E;
ram[9142] = 8'h43;
ram[9143] = 8'hB7;
ram[9144] = 8'h40;
ram[9145] = 8'h9E;
ram[9146] = 8'h86;
ram[9147] = 8'h9F;
ram[9148] = 8'h43;
ram[9149] = 8'hB7;
ram[9150] = 8'h40;
ram[9151] = 8'h9F;
ram[9152] = 8'h86;
ram[9153] = 8'hA0;
ram[9154] = 8'h43;
ram[9155] = 8'hB7;
ram[9156] = 8'h40;
ram[9157] = 8'hA0;
ram[9158] = 8'h86;
ram[9159] = 8'hA1;
ram[9160] = 8'h43;
ram[9161] = 8'hB7;
ram[9162] = 8'h40;
ram[9163] = 8'hA1;
ram[9164] = 8'h86;
ram[9165] = 8'hA2;
ram[9166] = 8'h43;
ram[9167] = 8'hB7;
ram[9168] = 8'h40;
ram[9169] = 8'hA2;
ram[9170] = 8'h86;
ram[9171] = 8'hA3;
ram[9172] = 8'h43;
ram[9173] = 8'hB7;
ram[9174] = 8'h40;
ram[9175] = 8'hA3;
ram[9176] = 8'h86;
ram[9177] = 8'hA4;
ram[9178] = 8'h43;
ram[9179] = 8'hB7;
ram[9180] = 8'h40;
ram[9181] = 8'hA4;
ram[9182] = 8'h86;
ram[9183] = 8'hA5;
ram[9184] = 8'h43;
ram[9185] = 8'hB7;
ram[9186] = 8'h40;
ram[9187] = 8'hA5;
ram[9188] = 8'h86;
ram[9189] = 8'hA6;
ram[9190] = 8'h43;
ram[9191] = 8'hB7;
ram[9192] = 8'h40;
ram[9193] = 8'hA6;
ram[9194] = 8'h86;
ram[9195] = 8'hA7;
ram[9196] = 8'h43;
ram[9197] = 8'hB7;
ram[9198] = 8'h40;
ram[9199] = 8'hA7;
ram[9200] = 8'h86;
ram[9201] = 8'hA8;
ram[9202] = 8'h43;
ram[9203] = 8'hB7;
ram[9204] = 8'h40;
ram[9205] = 8'hA8;
ram[9206] = 8'h86;
ram[9207] = 8'hA9;
ram[9208] = 8'h43;
ram[9209] = 8'hB7;
ram[9210] = 8'h40;
ram[9211] = 8'hA9;
ram[9212] = 8'h86;
ram[9213] = 8'hAA;
ram[9214] = 8'h43;
ram[9215] = 8'hB7;
ram[9216] = 8'h40;
ram[9217] = 8'hAA;
ram[9218] = 8'h86;
ram[9219] = 8'hAB;
ram[9220] = 8'h43;
ram[9221] = 8'hB7;
ram[9222] = 8'h40;
ram[9223] = 8'hAB;
ram[9224] = 8'h86;
ram[9225] = 8'hAC;
ram[9226] = 8'h43;
ram[9227] = 8'hB7;
ram[9228] = 8'h40;
ram[9229] = 8'hAC;
ram[9230] = 8'h86;
ram[9231] = 8'hAD;
ram[9232] = 8'h43;
ram[9233] = 8'hB7;
ram[9234] = 8'h40;
ram[9235] = 8'hAD;
ram[9236] = 8'h86;
ram[9237] = 8'hAE;
ram[9238] = 8'h43;
ram[9239] = 8'hB7;
ram[9240] = 8'h40;
ram[9241] = 8'hAE;
ram[9242] = 8'h86;
ram[9243] = 8'hAF;
ram[9244] = 8'h43;
ram[9245] = 8'hB7;
ram[9246] = 8'h40;
ram[9247] = 8'hAF;
ram[9248] = 8'h86;
ram[9249] = 8'hB0;
ram[9250] = 8'h43;
ram[9251] = 8'hB7;
ram[9252] = 8'h40;
ram[9253] = 8'hB0;
ram[9254] = 8'h86;
ram[9255] = 8'hB1;
ram[9256] = 8'h43;
ram[9257] = 8'hB7;
ram[9258] = 8'h40;
ram[9259] = 8'hB1;
ram[9260] = 8'h86;
ram[9261] = 8'hB2;
ram[9262] = 8'h43;
ram[9263] = 8'hB7;
ram[9264] = 8'h40;
ram[9265] = 8'hB2;
ram[9266] = 8'h86;
ram[9267] = 8'hB3;
ram[9268] = 8'h43;
ram[9269] = 8'hB7;
ram[9270] = 8'h40;
ram[9271] = 8'hB3;
ram[9272] = 8'h86;
ram[9273] = 8'hB4;
ram[9274] = 8'h43;
ram[9275] = 8'hB7;
ram[9276] = 8'h40;
ram[9277] = 8'hB4;
ram[9278] = 8'h86;
ram[9279] = 8'hB5;
ram[9280] = 8'h43;
ram[9281] = 8'hB7;
ram[9282] = 8'h40;
ram[9283] = 8'hB5;
ram[9284] = 8'h86;
ram[9285] = 8'hB6;
ram[9286] = 8'h43;
ram[9287] = 8'hB7;
ram[9288] = 8'h40;
ram[9289] = 8'hB6;
ram[9290] = 8'h86;
ram[9291] = 8'hB7;
ram[9292] = 8'h43;
ram[9293] = 8'hB7;
ram[9294] = 8'h40;
ram[9295] = 8'hB7;
ram[9296] = 8'h86;
ram[9297] = 8'hB8;
ram[9298] = 8'h43;
ram[9299] = 8'hB7;
ram[9300] = 8'h40;
ram[9301] = 8'hB8;
ram[9302] = 8'h86;
ram[9303] = 8'hB9;
ram[9304] = 8'h43;
ram[9305] = 8'hB7;
ram[9306] = 8'h40;
ram[9307] = 8'hB9;
ram[9308] = 8'h86;
ram[9309] = 8'hBA;
ram[9310] = 8'h43;
ram[9311] = 8'hB7;
ram[9312] = 8'h40;
ram[9313] = 8'hBA;
ram[9314] = 8'h86;
ram[9315] = 8'hBB;
ram[9316] = 8'h43;
ram[9317] = 8'hB7;
ram[9318] = 8'h40;
ram[9319] = 8'hBB;
ram[9320] = 8'h86;
ram[9321] = 8'hBC;
ram[9322] = 8'h43;
ram[9323] = 8'hB7;
ram[9324] = 8'h40;
ram[9325] = 8'hBC;
ram[9326] = 8'h86;
ram[9327] = 8'hBD;
ram[9328] = 8'h43;
ram[9329] = 8'hB7;
ram[9330] = 8'h40;
ram[9331] = 8'hBD;
ram[9332] = 8'h86;
ram[9333] = 8'hBE;
ram[9334] = 8'h43;
ram[9335] = 8'hB7;
ram[9336] = 8'h40;
ram[9337] = 8'hBE;
ram[9338] = 8'h86;
ram[9339] = 8'hBF;
ram[9340] = 8'h43;
ram[9341] = 8'hB7;
ram[9342] = 8'h40;
ram[9343] = 8'hBF;
ram[9344] = 8'h86;
ram[9345] = 8'hC0;
ram[9346] = 8'h43;
ram[9347] = 8'hB7;
ram[9348] = 8'h40;
ram[9349] = 8'hC0;
ram[9350] = 8'h86;
ram[9351] = 8'hC1;
ram[9352] = 8'h43;
ram[9353] = 8'hB7;
ram[9354] = 8'h40;
ram[9355] = 8'hC1;
ram[9356] = 8'h86;
ram[9357] = 8'hC2;
ram[9358] = 8'h43;
ram[9359] = 8'hB7;
ram[9360] = 8'h40;
ram[9361] = 8'hC2;
ram[9362] = 8'h86;
ram[9363] = 8'hC3;
ram[9364] = 8'h43;
ram[9365] = 8'hB7;
ram[9366] = 8'h40;
ram[9367] = 8'hC3;
ram[9368] = 8'h86;
ram[9369] = 8'hC4;
ram[9370] = 8'h43;
ram[9371] = 8'hB7;
ram[9372] = 8'h40;
ram[9373] = 8'hC4;
ram[9374] = 8'h86;
ram[9375] = 8'hC5;
ram[9376] = 8'h43;
ram[9377] = 8'hB7;
ram[9378] = 8'h40;
ram[9379] = 8'hC5;
ram[9380] = 8'h86;
ram[9381] = 8'hC6;
ram[9382] = 8'h43;
ram[9383] = 8'hB7;
ram[9384] = 8'h40;
ram[9385] = 8'hC6;
ram[9386] = 8'h86;
ram[9387] = 8'hC7;
ram[9388] = 8'h43;
ram[9389] = 8'hB7;
ram[9390] = 8'h40;
ram[9391] = 8'hC7;
ram[9392] = 8'h86;
ram[9393] = 8'hC8;
ram[9394] = 8'h43;
ram[9395] = 8'hB7;
ram[9396] = 8'h40;
ram[9397] = 8'hC8;
ram[9398] = 8'h86;
ram[9399] = 8'hC9;
ram[9400] = 8'h43;
ram[9401] = 8'hB7;
ram[9402] = 8'h40;
ram[9403] = 8'hC9;
ram[9404] = 8'h86;
ram[9405] = 8'hCA;
ram[9406] = 8'h43;
ram[9407] = 8'hB7;
ram[9408] = 8'h40;
ram[9409] = 8'hCA;
ram[9410] = 8'h86;
ram[9411] = 8'hCB;
ram[9412] = 8'h43;
ram[9413] = 8'hB7;
ram[9414] = 8'h40;
ram[9415] = 8'hCB;
ram[9416] = 8'h86;
ram[9417] = 8'hCC;
ram[9418] = 8'h43;
ram[9419] = 8'hB7;
ram[9420] = 8'h40;
ram[9421] = 8'hCC;
ram[9422] = 8'h86;
ram[9423] = 8'hCD;
ram[9424] = 8'h43;
ram[9425] = 8'hB7;
ram[9426] = 8'h40;
ram[9427] = 8'hCD;
ram[9428] = 8'h86;
ram[9429] = 8'hCE;
ram[9430] = 8'h43;
ram[9431] = 8'hB7;
ram[9432] = 8'h40;
ram[9433] = 8'hCE;
ram[9434] = 8'h86;
ram[9435] = 8'hCF;
ram[9436] = 8'h43;
ram[9437] = 8'hB7;
ram[9438] = 8'h40;
ram[9439] = 8'hCF;
ram[9440] = 8'h86;
ram[9441] = 8'hD0;
ram[9442] = 8'h43;
ram[9443] = 8'hB7;
ram[9444] = 8'h40;
ram[9445] = 8'hD0;
ram[9446] = 8'h86;
ram[9447] = 8'hD1;
ram[9448] = 8'h43;
ram[9449] = 8'hB7;
ram[9450] = 8'h40;
ram[9451] = 8'hD1;
ram[9452] = 8'h86;
ram[9453] = 8'hD2;
ram[9454] = 8'h43;
ram[9455] = 8'hB7;
ram[9456] = 8'h40;
ram[9457] = 8'hD2;
ram[9458] = 8'h86;
ram[9459] = 8'hD3;
ram[9460] = 8'h43;
ram[9461] = 8'hB7;
ram[9462] = 8'h40;
ram[9463] = 8'hD3;
ram[9464] = 8'h86;
ram[9465] = 8'hD4;
ram[9466] = 8'h43;
ram[9467] = 8'hB7;
ram[9468] = 8'h40;
ram[9469] = 8'hD4;
ram[9470] = 8'h86;
ram[9471] = 8'hD5;
ram[9472] = 8'h43;
ram[9473] = 8'hB7;
ram[9474] = 8'h40;
ram[9475] = 8'hD5;
ram[9476] = 8'h86;
ram[9477] = 8'hD6;
ram[9478] = 8'h43;
ram[9479] = 8'hB7;
ram[9480] = 8'h40;
ram[9481] = 8'hD6;
ram[9482] = 8'h86;
ram[9483] = 8'hD7;
ram[9484] = 8'h43;
ram[9485] = 8'hB7;
ram[9486] = 8'h40;
ram[9487] = 8'hD7;
ram[9488] = 8'h86;
ram[9489] = 8'hD8;
ram[9490] = 8'h43;
ram[9491] = 8'hB7;
ram[9492] = 8'h40;
ram[9493] = 8'hD8;
ram[9494] = 8'h86;
ram[9495] = 8'hD9;
ram[9496] = 8'h43;
ram[9497] = 8'hB7;
ram[9498] = 8'h40;
ram[9499] = 8'hD9;
ram[9500] = 8'h86;
ram[9501] = 8'hDA;
ram[9502] = 8'h43;
ram[9503] = 8'hB7;
ram[9504] = 8'h40;
ram[9505] = 8'hDA;
ram[9506] = 8'h86;
ram[9507] = 8'hDB;
ram[9508] = 8'h43;
ram[9509] = 8'hB7;
ram[9510] = 8'h40;
ram[9511] = 8'hDB;
ram[9512] = 8'h86;
ram[9513] = 8'hDC;
ram[9514] = 8'h43;
ram[9515] = 8'hB7;
ram[9516] = 8'h40;
ram[9517] = 8'hDC;
ram[9518] = 8'h86;
ram[9519] = 8'hDD;
ram[9520] = 8'h43;
ram[9521] = 8'hB7;
ram[9522] = 8'h40;
ram[9523] = 8'hDD;
ram[9524] = 8'h86;
ram[9525] = 8'hDE;
ram[9526] = 8'h43;
ram[9527] = 8'hB7;
ram[9528] = 8'h40;
ram[9529] = 8'hDE;
ram[9530] = 8'h86;
ram[9531] = 8'hDF;
ram[9532] = 8'h43;
ram[9533] = 8'hB7;
ram[9534] = 8'h40;
ram[9535] = 8'hDF;
ram[9536] = 8'h86;
ram[9537] = 8'hE0;
ram[9538] = 8'h43;
ram[9539] = 8'hB7;
ram[9540] = 8'h40;
ram[9541] = 8'hE0;
ram[9542] = 8'h86;
ram[9543] = 8'hE1;
ram[9544] = 8'h43;
ram[9545] = 8'hB7;
ram[9546] = 8'h40;
ram[9547] = 8'hE1;
ram[9548] = 8'h86;
ram[9549] = 8'hE2;
ram[9550] = 8'h43;
ram[9551] = 8'hB7;
ram[9552] = 8'h40;
ram[9553] = 8'hE2;
ram[9554] = 8'h86;
ram[9555] = 8'hE3;
ram[9556] = 8'h43;
ram[9557] = 8'hB7;
ram[9558] = 8'h40;
ram[9559] = 8'hE3;
ram[9560] = 8'h86;
ram[9561] = 8'hE4;
ram[9562] = 8'h43;
ram[9563] = 8'hB7;
ram[9564] = 8'h40;
ram[9565] = 8'hE4;
ram[9566] = 8'h86;
ram[9567] = 8'hE5;
ram[9568] = 8'h43;
ram[9569] = 8'hB7;
ram[9570] = 8'h40;
ram[9571] = 8'hE5;
ram[9572] = 8'h86;
ram[9573] = 8'hE6;
ram[9574] = 8'h43;
ram[9575] = 8'hB7;
ram[9576] = 8'h40;
ram[9577] = 8'hE6;
ram[9578] = 8'h86;
ram[9579] = 8'hE7;
ram[9580] = 8'h43;
ram[9581] = 8'hB7;
ram[9582] = 8'h40;
ram[9583] = 8'hE7;
ram[9584] = 8'h86;
ram[9585] = 8'hE8;
ram[9586] = 8'h43;
ram[9587] = 8'hB7;
ram[9588] = 8'h40;
ram[9589] = 8'hE8;
ram[9590] = 8'h86;
ram[9591] = 8'hE9;
ram[9592] = 8'h43;
ram[9593] = 8'hB7;
ram[9594] = 8'h40;
ram[9595] = 8'hE9;
ram[9596] = 8'h86;
ram[9597] = 8'hEA;
ram[9598] = 8'h43;
ram[9599] = 8'hB7;
ram[9600] = 8'h40;
ram[9601] = 8'hEA;
ram[9602] = 8'h86;
ram[9603] = 8'hEB;
ram[9604] = 8'h43;
ram[9605] = 8'hB7;
ram[9606] = 8'h40;
ram[9607] = 8'hEB;
ram[9608] = 8'h86;
ram[9609] = 8'hEC;
ram[9610] = 8'h43;
ram[9611] = 8'hB7;
ram[9612] = 8'h40;
ram[9613] = 8'hEC;
ram[9614] = 8'h86;
ram[9615] = 8'hED;
ram[9616] = 8'h43;
ram[9617] = 8'hB7;
ram[9618] = 8'h40;
ram[9619] = 8'hED;
ram[9620] = 8'h86;
ram[9621] = 8'hEE;
ram[9622] = 8'h43;
ram[9623] = 8'hB7;
ram[9624] = 8'h40;
ram[9625] = 8'hEE;
ram[9626] = 8'h86;
ram[9627] = 8'hEF;
ram[9628] = 8'h43;
ram[9629] = 8'hB7;
ram[9630] = 8'h40;
ram[9631] = 8'hEF;
ram[9632] = 8'h86;
ram[9633] = 8'hF0;
ram[9634] = 8'h43;
ram[9635] = 8'hB7;
ram[9636] = 8'h40;
ram[9637] = 8'hF0;
ram[9638] = 8'h86;
ram[9639] = 8'hF1;
ram[9640] = 8'h43;
ram[9641] = 8'hB7;
ram[9642] = 8'h40;
ram[9643] = 8'hF1;
ram[9644] = 8'h86;
ram[9645] = 8'hF2;
ram[9646] = 8'h43;
ram[9647] = 8'hB7;
ram[9648] = 8'h40;
ram[9649] = 8'hF2;
ram[9650] = 8'h86;
ram[9651] = 8'hF3;
ram[9652] = 8'h43;
ram[9653] = 8'hB7;
ram[9654] = 8'h40;
ram[9655] = 8'hF3;
ram[9656] = 8'h86;
ram[9657] = 8'hF4;
ram[9658] = 8'h43;
ram[9659] = 8'hB7;
ram[9660] = 8'h40;
ram[9661] = 8'hF4;
ram[9662] = 8'h86;
ram[9663] = 8'hF5;
ram[9664] = 8'h43;
ram[9665] = 8'hB7;
ram[9666] = 8'h40;
ram[9667] = 8'hF5;
ram[9668] = 8'h86;
ram[9669] = 8'hF6;
ram[9670] = 8'h43;
ram[9671] = 8'hB7;
ram[9672] = 8'h40;
ram[9673] = 8'hF6;
ram[9674] = 8'h86;
ram[9675] = 8'hF7;
ram[9676] = 8'h43;
ram[9677] = 8'hB7;
ram[9678] = 8'h40;
ram[9679] = 8'hF7;
ram[9680] = 8'h86;
ram[9681] = 8'hF8;
ram[9682] = 8'h43;
ram[9683] = 8'hB7;
ram[9684] = 8'h40;
ram[9685] = 8'hF8;
ram[9686] = 8'h86;
ram[9687] = 8'hF9;
ram[9688] = 8'h43;
ram[9689] = 8'hB7;
ram[9690] = 8'h40;
ram[9691] = 8'hF9;
ram[9692] = 8'h86;
ram[9693] = 8'hFA;
ram[9694] = 8'h43;
ram[9695] = 8'hB7;
ram[9696] = 8'h40;
ram[9697] = 8'hFA;
ram[9698] = 8'h86;
ram[9699] = 8'hFB;
ram[9700] = 8'h43;
ram[9701] = 8'hB7;
ram[9702] = 8'h40;
ram[9703] = 8'hFB;
ram[9704] = 8'h86;
ram[9705] = 8'hFC;
ram[9706] = 8'h43;
ram[9707] = 8'hB7;
ram[9708] = 8'h40;
ram[9709] = 8'hFC;
ram[9710] = 8'h86;
ram[9711] = 8'hFD;
ram[9712] = 8'h43;
ram[9713] = 8'hB7;
ram[9714] = 8'h40;
ram[9715] = 8'hFD;
ram[9716] = 8'h86;
ram[9717] = 8'hFE;
ram[9718] = 8'h43;
ram[9719] = 8'hB7;
ram[9720] = 8'h40;
ram[9721] = 8'hFE;
ram[9722] = 8'h86;
ram[9723] = 8'hFF;
ram[9724] = 8'h43;
ram[9725] = 8'hB7;
ram[9726] = 8'h40;
ram[9727] = 8'hFF;
ram[9728] = 8'h7E;
ram[9729] = 8'h26;
ram[9730] = 8'h00;
ram[65534] = 8'h20;
ram[65535] = 8'h00;


	end
	
	always @(rw or data_in)
	begin 
		ram[address] = (rw) ? ram[address] : data_in;
	end
	
	assign data_out = (rw) ? ram[address] : 8'bZZZZZZZZ;
	
endmodule

module hc11_test;
	
	reg reset;
	reg E;
	wire rw_w;
	wire [15:0] address_w;
	wire [7:0] data_w;
	wire [7:0] write_data_w;
	
	// Instantiate the microcontroller core and RAM and connect them together.
  	hc11cpu cpu1 (E, 1'b0, reset, 4'b0000, 1'b0,,,, rw_w, address_w, data_w, write_data_w,,,,,,,,);
	int_ram ram1 (E, rw_w, address_w, write_data_w, data_w);

	integer i;
	
  	logic [7:0] value;
	logic [7:0] expected_value;
    logic [7:0] index;
	
	initial
	begin	
		reset = 1'b0;
		E = 1'b0;
		
		// Reset the device.
		#5 reset = 1'b1;
		#5 reset = 1'b0;
			
		// Run the program for a finite amount of time.
		for (i = 0; i < 80000; i = i + 1)
		begin		
			#5 E = ~E;
			#5 E = ~E;
		end
		
		// Check the results of the program in RAM.
        
      	index = 0;
      
      	repeat (`MAX_INDEX)
		begin          
        
          // Check COMA starting at address $4000.
          value = ram1.ram[16'h4000 + index];
          expected_value = ~index;
          
          if (expected_value != value)
            $display ("Error in instruction LDAA or STAA. Value = %b, expected value = %b.", value, expected_value);
		
          // Complete the checks for remaining instructions.
          value = ram1.ram[16'h4100 + index];
          expected_value = ~index;
          
          if (expected_value != value)
            $display ("Error in instruction COMA. Value = %b, expected value = %b.", value, expected_value);
          
                    
          index++;
          
        end	
	end		
endmodule
